library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.tank_const.all;
use work.game_library.all;

entity tb_tank_control is
end tb_tank_control;

architecture testbench of tb_tank_control is
    -- Signals for the tank_control ports
    signal clk              : std_logic := '0';
    signal rst_n            : std_logic := '0';
    signal we               : std_logic := '0';
    signal tank_curr_pos_in : position := (0, 0);
    signal tank_next_pos_out: position;
    signal tank_display     : std_logic;
    signal tank_speed_in    : std_logic_vector(2 downto 0) := "001"; -- Speed = 1

    -- Testbench clock period
    constant clk_period : time := 10 ns;

begin

    -- Instantiate the tank_control module
    uut: entity work.tank_control
        port map(
            clk              => clk,
            rst_n            => rst_n,
            we               => we,
            tank_curr_pos_in => tank_curr_pos_in,
            tank_next_pos_out => tank_next_pos_out,
            tank_display     => tank_display,
            tank_speed_in    => tank_speed_in
        );

    -- Clock process
    clk_process: process
    begin
        while true loop
            clk <= '0';
            wait for clk_period / 2;
            clk <= '1';
            wait for clk_period / 2;
        end loop;
    end process;

    -- Testbench stimulus process
    stimulus_process: process
    begin
        -- Test Reset
        rst_n <= '1';
        wait for 2 * clk_period;
        rst_n <= '0';
        wait for clk_period;
		  --rst_n <= '0';
		  --wait for clk_period;

        -- Test Start State -> Move Right
        we <= '1';
        wait for 5 * clk_period; -- Allow time for transitions

        -- Test Move Right -> Move Left
        tank_curr_pos_in(0) <= 639 - TANK_WIDTH; -- Near right boundary
        wait for 2 * clk_period;
		  tank_curr_pos_in(0) <= 640 - TANK_WIDTH; -- Near right boundary
        wait for 2 * clk_period;

        -- Test Move Left -> Move Right
        tank_curr_pos_in(0) <= 1; -- Near left boundary
        wait for 2 * clk_period;
		  tank_curr_pos_in(0) <= 0; -- Near left boundary
        wait for 2 * clk_period;

        -- Test Die State
        we <= '0'; -- Simulate a condition to enter "die"
        wait for clk_period;
        tank_curr_pos_in(0) <= 0; -- Trigger die state
        wait for 5 * clk_period;

        -- Test Win State
        rst_n <= '0';
        wait for 2 * clk_period;
        rst_n <= '1';
        we <= '1';
        tank_curr_pos_in(0) <= 0; -- Reset to start state
        wait for clk_period;
        -- Add your win state condition here
        wait for 5 * clk_period;

        -- Test Done State
        -- Add appropriate conditions to simulate entering 'done'

        -- Finish simulation
        wait;
    end process;

end architecture testbench;
