library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.tank_const.all;
use work.game_library.all;

entity collision is
	port(
		clk, rst_n, we  : in std_logic;
		
		tank_pos_in : in position;
		bullet_pos_in      : in position;
		bullet_fired_in    : in std_logic;
		collsion_hit       : out std_logic;
		direction          : in std_logic
		--dead               : out std_logic;
		);
end entity collision;

architecture fsm of collision is

	-- Define the states, including 'done'
	type state_type is (start, check_hit, hit, win, done);
	signal current_state, next_state : state_type;

begin

	-- Asynchronous Reset and Synchronous State Update
	process(clk, rst_n)
		begin
			if rst_n = '1' then
				current_state <= start;
			elsif (rising_edge(clk)) then
				current_state <= next_state;
			end if;
	end process;
	
	-- Next State and Output Logic
	process(current_state, we, bullet_pos_in, bullet_fired_in, direction, tank_pos_in)
		--variable new_pos : position;
		--variable new_state : state_type;
	begin
		-- Default assignments to avoid latches
		next_state <= current_state;
		--collsion_hit <= ;
		--bullet_disp <= '0';
		
		case current_state is
		
			when start =>
				next_state <= check_hit;
				
				
			when check_hit =>
--				if we = '1' then
--					if direction = '0' then
--						bullet_pos_out(1) <= bullet_pos_in(1) - speed;
--						bullet_pos_out(0) <= bullet_pos_in(0);
--					else
--						bullet_pos_out(1) <= bullet_pos_in(1) + speed;
--						bullet_pos_out(0) <= bullet_pos_in(0);
--					end if;
--				end if;
				if (((tank_pos_in(1) > tank_1_pos_in(1) - TANK_GUNH) 
					   and (tank_pos_in(1) - BULLET_H < tank_1_pos_in(1) + TANK_HEIGHT) 
					   and (tank_pos_in(0) - BULLET_W/2 < tank_1_pos_in(0) + TANK_WIDTH) 
					   and (tank_pos_in(0) + BULLET_W/2 > tank_1_pos_in(0))
					   and bul_2_hit = '0')) then
					next_state <= hit_boundary;
				else
					next_state <= move_bullet;
				end if;
				bullet_fired_out <= '1';
			
			when hit_boundary =>
				next_state <= start;
			   bullet_disp <= '0'; -- Turn off display	
				bullet_fired_out <= '0';
				bullet_pos_out(0) <= -1000;
				bullet_pos_out(1) <= -1000;
			
			when die =>
				bullet_disp <= '0'; -- Turn off display
				next_state <= done;
				bullet_pos_out(0) <= -1000;
				bullet_pos_out(1) <= -1000;
				bullet_fired_out <= '0';
			
			when win =>
				bullet_disp <= '1'; -- Keep display ON
				next_state <= done;
				bullet_pos_out <= bullet_pos_in;
				bullet_fired_out <= '1';
			
			when done =>
				-- Maintain the current state values explicitly
				next_state <= done;
				bullet_pos_out(0) <= -1000;
				bullet_pos_out(1) <= -1000;
				bullet_fired_out <= '0';
			
			when others =>
				-- Explicitly assign defaults in case of unexpected state
				next_state <= start;
				bullet_disp <= '1';
				bullet_pos_out(0) <= 300;
				bullet_pos_out(1) <= 300;
				bullet_fired_out <= '0';
				
			end case;
	end process;

end architecture fsm;