library IEEE;
use IEEE.std_logic_1164.all;

package game_library is
	type position is array(0 to 1) of integer;
	
end package game_library;

package body game_library is
end package body game_library;