

entity tankgame is

end entity tankgame;